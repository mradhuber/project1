module ps4(	
	input		 [3:0] req,
	input		  	   en,
	output logic [3:0] gnt
);

// using if statements